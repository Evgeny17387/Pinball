module tb

endmodule
