package score;

    localparam TOP_SCORES_NUM = 3;

endpackage
