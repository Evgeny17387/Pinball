
const int xFrameSize = 635;
const int yFrameSize = 475;
