
parameter logic [7:0] BUMPER_COLOR = 8'b01010111;
