parameter logic [10:0] LIFE_TOP_LEFT_X = 30;
parameter logic [10:0] LIFE_TOP_LEFT_Y = 5;

localparam LIFE_SPACE = 40;

parameter logic [10:0] SCORE_TOP_LEFT_X = 170;
parameter logic [10:0] SCORE_TOP_LEFT_Y = 5;

parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_X = 220;
parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_Y = 5;
