import defines::COLOR_TRANSPARENT, defines::COLOR_YELLOW;

module score_bitmap(	
	input	logic			clk,
	input	logic			resetN,
	input 	logic	[10:0] 	offsetX,
	input 	logic	[10:0] 	offsetY,
	input	logic			insideRectangle,
	output	logic			drawStar,
	output	logic	[7:0] 	RGBStar
);

`ifdef PICTURES
logic[0:31][0:31] object_colors = {
	32'b11111111111111111111111111111111,
	32'b11111111111111101111111111111111,
	32'b11111111111111100111111111111111,
	32'b11111111111111000111111111111111,
	32'b11111111111111000011111111111111,
	32'b11111111111110000011111111111111,
	32'b11111111111110000001111111111111,
	32'b11111111111100000001111111111111,
	32'b11111111111100000000111111111111,
	32'b11111111111000000000111111111111,
	32'b11111111111000000000011111111111,
	32'b11111000000000000000000000011111,
	32'b00000000000000000000000000000000,
	32'b10000000000000000000000000000001,
	32'b11000000000000000000000000000011,
	32'b11100000000000000000000000000111,
	32'b11110000000000000000000000001111,
	32'b11111000000000000000000000011111,
	32'b11111100000000000000000000111111,
	32'b11111110000000000000000001111111,
	32'b11111111000000000000000011111111,
	32'b11111111000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000001111111,
	32'b11111110000000000000000001111111,
	32'b11111110000000000000000001111111,
	32'b11111110000000011000000001111111,
	32'b11111110000001111110000001111111,
	32'b11111100000111111111100001111111,
	32'b11111100011111111111111000111111,
	32'b11111101111111111111111110111111,
	32'b11111111111111111111111111111111};
`endif

always_ff@(posedge clk or negedge resetN)
begin

	if (!resetN) begin
		RGBStar <= 8'h00;
	end

	else begin

		RGBStar <= COLOR_TRANSPARENT;

		if (insideRectangle == 1'b1) begin

`ifdef PICTURES
			RGBStar <= (object_colors[offsetY][offsetX] ==  0) ? COLOR_YELLOW : COLOR_TRANSPARENT;
`else
			RGBStar <= COLOR_YELLOW;
`endif

		end
	end

end

assign drawStar = (RGBStar != COLOR_TRANSPARENT) ? 1'b1 : 1'b0;

endmodule
