localparam WORD_WELCOME_TOP_LEFT_X = 150;
localparam WORD_WELCOME_TOP_LEFT_Y = 50;
localparam WORD_WELCOME_SIZE = 8;
localparam int WORD_WELCOME_LETTERS[WORD_WELCOME_SIZE-1:0] = '{4, 12, 14, 2, 11, 11, 4, 22};

localparam WORD_WELCOME_2_TOP_LEFT_X = 1;
localparam WORD_WELCOME_2_TOP_LEFT_Y = 150;
localparam WORD_WELCOME_2_SIZE = 13;
localparam int WORD_WELCOME_2_LETTERS[WORD_WELCOME_2_SIZE-1:0] = '{27, 4, 15, 24, 19, 26, 17, 4, 15, 15, 8, 11, 5};

localparam WORD_WELCOME_3_TOP_LEFT_X = 100;
localparam WORD_WELCOME_3_TOP_LEFT_Y = 250;
localparam WORD_WELCOME_3_SIZE = 6;
localparam int WORD_WELCOME_3_LETTERS[WORD_WELCOME_3_SIZE-1:0] = '{4, 11, 6, 13, 8, 18};

localparam WORD_WELCOME_4_TOP_LEFT_X = 400;
localparam WORD_WELCOME_4_TOP_LEFT_Y = 250;
localparam WORD_WELCOME_4_SIZE = 4;
localparam int WORD_WELCOME_4_LETTERS[WORD_WELCOME_4_SIZE-1:0] = '{11, 0, 20, 3};

localparam WORD_WELCOME_5_TOP_LEFT_X = 1;
localparam WORD_WELCOME_5_TOP_LEFT_Y = 350;
localparam WORD_WELCOME_5_SIZE = 10;
localparam int WORD_WELCOME_5_LETTERS[WORD_WELCOME_5_SIZE-1:0] = '{27, 3, 8, 26, 17, 4, 24, 0, 11, 15};

localparam SCREEN_WELCOME_PLAYER_ID_TOP_LEFT_X = 100;
localparam SCREEN_WELCOME_PLAYER_ID_TOP_LEFT_Y = 425;
