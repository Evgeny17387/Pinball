
parameter logic [10:0] SCORE_TOP_LEFT_X = 120;
parameter logic [10:0] SCORE_TOP_LEFT_Y = 5;
