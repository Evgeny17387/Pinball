
parameter logic [7:0] COLOR_TRANSPARENT = 8'b11111111;

parameter logic [7:0] COLOR_RED         = 8'b11000000;
parameter logic [7:0] COLOR_GREEN       = 8'b00111000;
parameter logic [7:0] COLOR_BLUE        = 8'b00000111;
parameter logic [7:0] COLOR_WHITE       = 8'b11111111;
parameter logic [7:0] COLOR_BLACK       = 8'b00000000;
parameter logic [7:0] COLOR_YELLOW      = 8'b11111000;
parameter logic [7:0] COLOR_BLUE_DARK   = 8'h11101101;
parameter logic [7:0] COLOR_PURPLE        = 8'b10110011;

parameter logic [7:0] COLOR_DEFAULT     = 8'b01011011;
