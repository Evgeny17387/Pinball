
const int FRAME_SIZE_X = 635;
const int FRAME_SIZE_Y = 475;

const int FIXED_POINT_MULTIPLIER = 64;
