
localparam LIFE_INIT = 3;
