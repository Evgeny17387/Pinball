
parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_X = 70;
parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_Y = 5;

parameter logic [10:0] LEVEL_LABEL_TOP_LEFT_X = 20;
parameter logic [10:0] LEVEL_LABEL_TOP_LEFT_Y = 5;

parameter logic [10:0] LEVEL_LABEL_WIDTH = 16;
parameter logic [10:0] LEVEL_LABEL_HEIGHT = 16;

parameter logic [7:0] LEVEL_LABEL_COLOR = 8'hAA;
