
typedef struct packed {
	logic signed [3:0] xxFactor;
	logic signed [3:0] xyFactor;
	logic signed [3:0] yyFactor;
	logic signed [3:0] yxFactor;
} COLLISION_FACTOR;
