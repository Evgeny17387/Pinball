
parameter logic [7:0] BUMPER_COLOR = COLOR_BLUE;
