
localparam SPRING_SPEED_DOWN = 50;
localparam SPRING_SPEED_UP = -100;

localparam SPRING_Y_MARGIN = 20;
