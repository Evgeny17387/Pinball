
localparam LETTER_SPACE = 40;
