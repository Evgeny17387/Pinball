
localparam LIFE_INIT = 2;
