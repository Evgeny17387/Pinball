
const int FIXED_POINT_MULTIPLIER = 64;
