
const int GRAVITY = 5;

parameter logic [7:0] BALL_COLOR = COLOR_BLUE_DARK;
