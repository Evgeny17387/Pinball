package defines;

    parameter int INITIAL_X = 280;
    parameter int INITIAL_Y = 185;

    parameter logic signed [10:0] SCORE_TOP_LEFT_X = 50;
    parameter logic signed [10:0] SCORE_TOP_LEFT_Y = 50;

    parameter logic signed [10:0] LEVEL_TOP_LEFT_X = 50;
    parameter logic signed [10:0] LEVEL_TOP_LEFT_Y = 100;

    parameter logic signed [10:0] LEVEL_STATUS_TOP_LEFT_X = 550;
    parameter logic signed [10:0] LEVEL_STATUS_TOP_LEFT_Y = 50;

endpackage
