
const int bracketOffset_h = 10;
const int bracketOffset_top = 50;
const int bracketOffset_bottom = 10;
