
localparam SPRING_SPEED_DOWN = 100;
localparam SPRING_SPEED_UP = -200;

localparam SPRING_Y_MARGIN = 20;
