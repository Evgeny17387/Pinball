
parameter logic [10:0]  NUMBER_WIDTH    = 16;
parameter logic [10:0]  NUMBER_HEIGHT   = 32;

parameter logic [10:0]  NUMBER_SPACE    = 20;
