
parameter logic [10:0] LIFE_NUMBER_TOP_LEFT_X = 170;
parameter logic [10:0] LIFE_NUMBER_TOP_LEFT_Y = 5;
