import defines::LIFE_WIDTH, defines::LIFE_HEIGHT;
import defines::COLOR_TRANSPARENT, defines::COLOR_RED;

module life_bitmap(
    input   logic	        clk,
    input	logic	        resetN,
    input   logic	[10:0]  offsetX,
    input   logic	[10:0]  offsetY,
    input	logic	        insideRectangle,
    output	logic	        drawLife,
    output	logic	[7:0]   RGBLife
);

logic[0:LIFE_HEIGHT-1][0:LIFE_WIDTH-1] object_colors = {
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000011111100000000111111000000,
	32'b00001111111111000011111111110000,
	32'b00011111111111100111111111111000,
	32'b00011111111111111111111111111000,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00111111111111111111111111111100,
	32'b00011111111111111111111111111000,
	32'b00011111111111111111111111111000,
	32'b00001111111111111111111111110000,
	32'b00001111111111111111111111100000,
	32'b00000111111111111111111111000000,
	32'b00000011111111111111111110000000,
	32'b00000000111111111111111100000000,
	32'b00000000011111111111111000000000,
	32'b00000000001111111111110000000000,
	32'b00000000000111111111100000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000001111110000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000000010000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
};

always_ff@(posedge clk or negedge resetN) 
begin 

	if(!resetN) begin 
		RGBLife <=	8'h00; 
	end 
	else begin 
		RGBLife <= COLOR_TRANSPARENT;

		if (insideRectangle == 1'b1)
		begin
			RGBLife <= (object_colors[offsetY][offsetX] ==  1) ? COLOR_RED : COLOR_TRANSPARENT;
		end

	end
end

assign drawLife = (RGBLife != COLOR_TRANSPARENT ) ? 1'b1 : 1'b0 ;

endmodule
