
parameter logic [7:0] TRAP_COLOR = COLOR_NEW;
