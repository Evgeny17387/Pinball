
localparam SPRING_SPEED_DOWN = 200;
localparam SPRING_SPEED_UP = -400;
