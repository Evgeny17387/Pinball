
parameter logic [7:0] FLIPPER_COLOR = COLOR_DEFAULT;
