
localparam LIFE_INIT = 1;
