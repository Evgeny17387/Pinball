// Life

parameter logic [10:0] LIFE_WIDTH = 32;
parameter logic [10:0] LIFE_HEIGHT = 32;

parameter logic [10:0] LIFE_TOP_LEFT_X = 30;
parameter logic [10:0] LIFE_TOP_LEFT_Y = 5;

localparam LIFE_SPACE = 40;

// Score

parameter logic [10:0] SCREEN_MAIN_SCORE_WIDTH = 32;
parameter logic [10:0] SCREEN_MAIN_SCORE_HEIGHT = 32;

parameter logic [10:0] SCREEN_MAIN_SCORE_TOP_LEFT_X = 170;
parameter logic [10:0] SCREEN_MAIN_SCORE_TOP_LEFT_Y = 5;

parameter logic [10:0] SCREEN_MAIN_SCORE_NUMBER_TOP_LEFT_X = 220;
parameter logic [10:0] SCREEN_MAIN_SCORE_NUMBER_TOP_LEFT_Y = 5;

// Level

parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_X = 300;
parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_Y = 5;

// Equation

parameter logic [10:0] SCREEN_MAIN_LUCK_SYMBOL_WIDTH = 32;
parameter logic [10:0] SCREEN_MAIN_LUCK_SYMBOL_HEIGHT = 32;

parameter logic [10:0] SCREEN_MAIN_LUCK_SYMBOL_TOP_LEFT_X = 450;
parameter logic [10:0] SCREEN_MAIN_LUCK_SYMBOL_TOP_LEFT_Y = 5;

parameter logic [10:0] SCREEN_MAIN_LUCK_NUMBER_TOP_LEFT_X = 500;
parameter logic [10:0] SCREEN_MAIN_LUCK_NUMBER_TOP_LEFT_Y = 5;

// Spring

parameter logic [10:0] SCREEN_MAIN_SPRING_WIDTH = 64;
parameter logic [10:0] SCREEN_MAIN_SPRING_HEIGHT = 220;

parameter logic [10:0] SCREEN_MAIN_SPRING_TOP_LEFT_X = 550;
parameter logic [10:0] SCREEN_MAIN_SPRING_TOP_LEFT_Y = 275;

// Ball

parameter int SCREEN_MAIN_BALL_INITIAL_X = 550;
parameter int SCREEN_MAIN_BALL_INITIAL_Y = 212;
