
localparam SPRING_SPEED_DOWN = 100;
localparam SPRING_SPEED_UP = -200;
