
localparam SPRING_SPEED = 5;

localparam SPRING_Y_MARGIN = 20;
