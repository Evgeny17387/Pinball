import defines::COLOR_TRANSPARENT, defines::COLOR_DEFAULT;
import defines::LETTER_HEIGHT, defines::LETTER_WIDTH;

module letter
#(parameter TOP_LEFT_X = 0, TOP_LEFT_Y = 0)
(
	input 	logic 			clk,
	input 	logic 			resetN,
	input 	logic	[10:0]	pixelX,
	input 	logic	[10:0]	pixelY,
	input	logic	[3:0] 	letter,
	output	logic			drawLetter,
	output	logic	[7:0]	RGBLetter
);

`ifdef PICTURES
bit [0:1] [0:LETTER_HEIGHT - 1] [0:LETTER_WIDTH - 1] letter_bitmap = {
// A - 0
{
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111
},
// B - 1
{
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000
}
};
`endif

logic insideLetter;

assign insideLetter = ((pixelX >= TOP_LEFT_X) && (pixelX < TOP_LEFT_X + LETTER_WIDTH) && (pixelY >= TOP_LEFT_Y) && (pixelY < TOP_LEFT_Y + LETTER_HEIGHT));

always_ff@(posedge clk or negedge resetN)
begin

	if(!resetN) begin

		drawLetter <= 1'b0;

	end
	else begin

		drawLetter <= 1'b0;

		if (insideLetter == 1'b1)

`ifdef PICTURES
			drawLetter <= (letter_bitmap[letter][pixelY - TOP_LEFT_Y][pixelX - TOP_LEFT_X]);
`else
			drawLetter <= 1'b1;
`endif

	end

end

assign RGBLetter = COLOR_DEFAULT;

endmodule 
