
localparam WORD_END_TOP_LEFT_X = 125;
localparam WORD_END_TOP_LEFT_Y = 100;
localparam WORD_END_SIZE = 9;
localparam int WORD_END_LETTERS[WORD_END_SIZE-1:0] = '{17, 4, 21, 14, 26, 4, 12, 0, 6};

localparam WORD_END_2_TOP_LEFT_X = 10;
localparam WORD_END_2_TOP_LEFT_Y = 300;
localparam WORD_END_2_SIZE = 14;
localparam int WORD_END_2_LETTERS[WORD_END_2_SIZE-1:0] = '{27, 18, 8, 26, 4, 17, 14, 2, 18, 26, 17, 20, 14, 24};

parameter logic [10:0] SCORE_NUMBER_TOP_LEFT_X = 10;
parameter logic [10:0] SCORE_NUMBER_TOP_LEFT_Y = 400;
