
const int GRAVITY = 2;
