package defines;

    parameter int INITIAL_X = 280;
    parameter int INITIAL_Y = 185;

endpackage
