
const int GRAVITY = 5;
