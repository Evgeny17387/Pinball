import defines::COLOR_TRANSPARENT, defines::COLOR_DEFAULT;
import defines::LETTER_HEIGHT, defines::LETTER_WIDTH;

module letter
(
	input 	logic 			clk,
	input 	logic 			resetN,
	input 	logic	[10:0]	offsetX,
	input 	logic	[10:0]	offsetY,
	input	logic	[3:0] 	letter,
	input 	logic 			drawLetter,
	output	logic			drawLetterBitMask,
	output	logic	[7:0]	RGBLetter
);

`ifdef PICTURES
// A - 0
// B - 1
bit [0:1] [0:LETTER_HEIGHT - 1] [0:LETTER_WIDTH - 1] letter_bitmap = {
// A - 0
{
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111,
	32'b11111110000000000000000011111111
},
// B - 1
{
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111100000000000000000001111111,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000,
	32'b11111111111111111111111111000000
}
};
`endif

always_ff@(posedge clk or negedge resetN)
begin

	if(!resetN) begin

		drawLetterBitMask <= 1'b0;

	end
	else begin

		drawLetterBitMask <= 1'b0;

		if (drawLetter == 1'b1)

`ifdef PICTURES
			drawLetterBitMask <= (letter_bitmap[letter][offsetY][offsetX]);
`else
			drawLetterBitMask <= 1'b1;
`endif

	end

end

assign RGBLetter = COLOR_DEFAULT;

endmodule 
