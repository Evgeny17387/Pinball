import defines::SCREEN_MAIN_LUCK_SYMBOL_WIDTH, defines::SCREEN_MAIN_LUCK_SYMBOL_HEIGHT;
import defines::COLOR_TRANSPARENT, defines::COLOR_GREEN;

module luck_bitmap(
    input   logic	        clk,
    input	logic	        resetN,
    input   logic	[10:0]  offsetX,
    input   logic	[10:0]  offsetY,
    input	logic	        insideRectangle,
    output	logic	        drawLuck,
    output	logic	[7:0]   RGBLuck
);

logic[0:SCREEN_MAIN_LUCK_SYMBOL_HEIGHT-1][0:SCREEN_MAIN_LUCK_SYMBOL_WIDTH-1] object_colors = {
	32'b00000000000000000000111111000000,
	32'b00000000000000000001111111100000,
	32'b00000111111110000011111111111000,
	32'b00000111111111000111111111111110,
	32'b01111111111111100111111111111111,
	32'b11111111111111110111111111111111,
	32'b11111111111111111111111111111110,
	32'b11111111111111111111111111111110,
	32'b11111111111111110111111111111100,
	32'b01111111111111110111111111111000,
	32'b00001111111111110111111111000000,
	32'b00000000000111111111000011000000,
	32'b00001111111111111111111111111000,
	32'b00011111111111111111111111111110,
	32'b00111111111111111111111111111111,
	32'b00111111111111110111111111111111,
	32'b01111111111111110111111111111111,
	32'b01111111111111110101111111111111,
	32'b01111111111111110101111111111110,
	32'b00111111111111110100111111111100,
	32'b00001111111111100100011111111100,
	32'b00001111111111001100001111111100,
	32'b00000111111110001000000001110000,
	32'b00000001111000001000000000000000,
	32'b00000000000000001000000000000000,
	32'b00000000000000001000000000000000,
	32'b00000000000000001000000000000000,
	32'b00000000000000011000000000000000,
	32'b00000000000000010000000000000000,
	32'b00000000000000010000000000000000,
	32'b00000000000000110000000000000000,
	32'b00000000000000100000000000000000
};

always_ff@(posedge clk or negedge resetN) 
begin 

	if(!resetN) begin 
		RGBLuck <=	8'h00; 
	end 
	else begin 
		RGBLuck <= COLOR_TRANSPARENT;

		if (insideRectangle == 1'b1)
		begin
			RGBLuck <= (object_colors[offsetY][offsetX] ==  1) ? COLOR_GREEN : COLOR_TRANSPARENT;
		end

	end
end

assign drawLuck = (RGBLuck != COLOR_TRANSPARENT ) ? 1'b1 : 1'b0 ;

endmodule
