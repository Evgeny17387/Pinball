
localparam logic [2:0]  COLOR_DARK              = 3'b111;
localparam logic [2:0]  COLOR_LIGHT             = 3'b000;

parameter logic [7:0]   COLOR_TRANSPARENT       = 8'hFF;
parameter logic [7:0] 	COLOR_DEFAULT 			= 8'h5b;

parameter logic [7:0] 	COLOR_WHITE 			= 8'hFF;
parameter logic [7:0] 	COLOR_RED 			    = 8'b11000000;
parameter logic [7:0] 	COLOR_YELLOW		    = 8'b11111000;
