
parameter logic [10:0] LETTER_WIDTH = 32;
parameter logic [10:0] LETTER_HEIGHT = 32;
