
parameter int INITIAL_Y_SPEED = 200;
