
parameter logic [7:0] COLOR_TRANSPARENT = 8'hFF;

parameter logic [7:0] COLOR_RED         = 8'b11000000;
parameter logic [7:0] COLOR_GREEN       = 8'b00111000;
parameter logic [7:0] COLOR_BLUE        = 8'b00000111;

parameter logic [7:0] COLOR_WHITE       = 8'hFF;
parameter logic [7:0] COLOR_YELLOW      = 8'b11111000;

parameter logic [7:0] COLOR_BLACK       = 8'h00;
parameter logic [7:0] COLOR_GRAY        = 8'h10010010;

parameter logic [7:0] COLOR_DEFAULT     = 8'h5b;
