
const int GRAVITY = 1;
