parameter logic [10:0] LIFE_TOP_LEFT_X = 170;
parameter logic [10:0] LIFE_TOP_LEFT_Y = 5;

localparam LIFE_SPACE = 40;
