
parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_X = 70;
parameter logic [10:0] LEVEL_NUMBER_TOP_LEFT_Y = 5;
