module tb_word

square #(.TOP_LEFT_X(250), .TOP_LEFT_Y(5)) square_inst(

);

initial begin
    #5 

end

endmodule
